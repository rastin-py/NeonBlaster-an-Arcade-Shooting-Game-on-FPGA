library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

package NeonBlaster_pkg is

type NumbersMap is array (0 to 15) of std_logic_vector(0 to 7);
type PlayerMap is array (0 to 34) of std_logic_vector(0 to 49);
type ShotsMap is array (0 to 7) of std_logic_vector(0 to 7);

--constant MAP_PLAYER : PlayerMap := (
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000000000000000000000000000000000000", -- 0
--    "00000000000000000011100000000111000000000000000000", -- 0
--    "00000000000000000110000000000001100000000000000000", -- 0
--    "00000000000000011100000000000000111000000000000000", -- 0
--    "00000000000001110000000000000000001110000000000000", -- 0
--    "00000000000011100000000000000000000111000000000000", --0 
--    "00000000001111000000000000000000000011100000000000", -- 0
--    "00000000011110000000000000000000000000111000000000", -- 0
--    "00000001111100000000000000000000000000001110000000", -- 0
--    "00000111110000000000000000000000000000001111100000", -- 0
--    "00001111100000000000000000000000000000000111110000", -- 0
--    "00011111100000000001000000000010000000000011111000", -- 0
--    "00011111100000000011100000000111000000000111111000", -- 0
--    "00111111110000000111110000001111100000001111111100", -- 0
--    "01111111111000001111111000011111110000011111111110", -- 0
--    "01111111111100011111111100111111111000111111111110", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "11111111111111111111111111111111111111111111111111", -- 0
--    "01111111111111111111111111111111111111111111111110", -- 0
--    "00111111111111111111111100111111111111111111111100", -- 0
--    "00001111111111111111111000011111111111111111110000", -- 0
--    "00000001111111111111100000000111111111111110000000", -- 0
--    "00000000011111111110000000000001111111111000000000", -- 0
--    "00000000000001111100000000000000111110000000000000", -- 0
--    "00000000000000111000000000000000011100000000000000" -- 0
--    );

constant MAP_PLAYER : PlayerMap := (
    "00000000000000000000111100001110000000000000000000", -- 0
    "00000000000000000111100000000111100000000000000000", -- 0
    "00000000000000111100000000000000111100000000000000", --0 
    "00000000000111110000000000000000001111100000000000", -- 0
    "00000000011111000000000000000000000011111000000000", -- 0
    "00000001111100000000000000000000000000111110000000", -- 0
    "00000011111000000000000000000000000000011111000000", -- 0
    "00001111110000000000000000000000000000001111110000", -- 0
    "00011111100000000001000000000010000000000111111000", -- 0
    "00111111100000000011100000000111000000000111111100", -- 0
    "01111111100000000111110000001111100000000111111110", -- 0
    "11111111110000001111111000011111110000001111111111", -- 0
    "11111111111000011111111100111111111000011111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "11111111111111111111111111111111111111111111111111", -- 0
    "01111111111111111111111111111111111111111111111110", -- 0
    "01111111111111111111111111111111111111111111111110", -- 0
    "00111111111111111111111111111111111111111111111100", -- 0
    "00011111111111111111111111111111111111111111111000", -- 0
    "00001111111111111111111111111111111111111111110000", -- 0
    "00000111111111111111111111111111111111111111100000", -- 0
    "00000011111111111111111111111111111111111111000000", -- 0
    "00000001111111111111100000000111111111111110000000", -- 0
    "00000000111111111110000000000001111111111100000000", -- 0
    "00000000011111111000000000000000011111111000000000", -- 0
    "00000000001111110000000000000000001111110000000000", -- 0
    "00000000000111100000000000000000000111100000000000", -- 0
    "00000000000011100000000000000000000111000000000000", -- 0
    "00000000000001110000000000000000001110000000000000",  
    "00000000000000011000000000000000011000000000000000", -- 
    "00000000000000000100000000000000100000000000000000" --  
    );
constant MAP_ZERO : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"11000110", -- 6 **   **
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000" -- f
		);
		
constant MAP_ONE : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"00011000", -- 2
		"00111000", -- 3
		"01111000", -- 4    **
		"00011000", -- 5   ***
		"00011000", -- 6  ****
		"00011000", -- 7    **
		"00011000", -- 8    **
		"00011000", -- 9    **
		"00011000", -- a    **
		"01111110", -- b    **
		"00000000", -- c    **
		"00000000", -- d  ******
		"00000000", -- e
		"00000000"  -- f
		);

constant MAP_TWO : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00001100", -- 5     **
		"00011000", -- 6    **
		"00110000", -- 7   **
		"01100000", -- 8  **
		"11000000", -- 9 **
		"11000110", -- a **   **
		"11111110", -- b *******
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
		);
		
constant MAP_THREE : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00111100", -- 6   ****
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
		);
		
constant MAP_FOUR : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"00001100", -- 2     **
		"00011100", -- 3    ***
		"00111100", -- 4   ****
		"01101100", -- 5  ** **
		"11001100", -- 6 **  **
		"11111110", -- 7 *******
		"00001100", -- 8     **
		"00001100", -- 9     **
		"00001100", -- a     **
		"00011110", -- b    ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
		);
		
constant MAP_FIVE : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000000", -- 3 **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
		);
		
constant MAP_SIX : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"00111000", -- 2   ***
		"01100000", -- 3  **
		"11000000", -- 4 **
		"11000000", -- 5 **
		"11111100", -- 6 ******
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000"  -- f
		);
		
constant MAP_SEVEN : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"11111110", -- 2 *******
		"11000110", -- 3 **   **
		"00000110", -- 4      **
		"00000110", -- 5      **
		"00001100", -- 6     **
		"00011000", -- 7    **
		"00110000", -- 8   **
		"00110000", -- 9   **
		"00110000", -- a   **
		"00110000", -- b   **
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000" -- f
		);
		
constant MAP_EIGHT : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111100", -- 6  *****
		"11000110", -- 7 **   **
		"11000110", -- 8 **   **
		"11000110", -- 9 **   **
		"11000110", -- a **   **
		"01111100", -- b  *****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000" -- f
		);
		
constant MAP_NINE : NumbersMap := (
		"00000000", -- 0
		"00000000", -- 1
		"01111100", -- 2  *****
		"11000110", -- 3 **   **
		"11000110", -- 4 **   **
		"11000110", -- 5 **   **
		"01111110", -- 6  ******
		"00000110", -- 7      **
		"00000110", -- 8      **
		"00000110", -- 9      **
		"00001100", -- a     **
		"01111000", -- b  ****
		"00000000", -- c
		"00000000", -- d
		"00000000", -- e
		"00000000" -- f
		);
		
constant MAP_SHOT : ShotsMap := (
		"00011000", -- 0
		"00111100", -- 1
		"01111110", -- 2
		"11111111", -- 3
		"11111111", -- 4    *
		"11111111", -- 5   ***
		"11111111", -- 6   ***
		"11111111" -- 7   
		);
type healthMapType is array (0 to 9) of NumbersMap;
constant HEALTH_MAP : healthMapType := (MAP_ZERO, MAP_ONE, MAP_TWO, MAP_THREE, MAP_FOUR, MAP_FIVE, MAP_SIX, MAP_SEVEN, MAP_EIGHT, MAP_NINE);
type EnemyType is record
  x_position        : integer;   -- X position of the enemy
  y_position        : integer;   -- Y position of the enemy
  x_speed           : integer;   -- X speed of the enemy
  y_speed           : integer;   -- Y speed of the enemy
  x_direction       : std_logic;   -- X direction of the enemy
  y_direction       : std_logic;   -- Y direction of the enemy
  gravity           : integer;   -- Gravity affecting the enemy
  color             : std_logic_vector(2 downto 0);   -- Color of the enemy
  is_alive          : std_logic;   -- Indicates whether the enemy is alive
  spawning          : std_logic;   -- Indicates whether the enemy is under attack
  health            : integer;   -- Health of the enemy
  initial_health    : integer;   -- Health of the enemy
end record;
type EnemyArrayType is array (natural range <>) of EnemyType;

type PlayerType is record
  x_position       : integer;
  y_position       : integer;
  is_alive         : std_logic;
  score            : integer;
end record;

type ShotType is record
  x_position      : integer;
  y_position      : integer;
  segment         : integer;
  iterator        : integer;
end record;

type BombType is record
  x_position      : integer;
  y_position      : integer;
  hit             : std_logic;
end record;
type BombArrayType is array (natural range <>) of BombType;

type GameStateType is (HOLD, STARTED, ENDED);
type GameType is record
  state      : GameStateType;
  timer           : integer;
  enemies_killed   : integer;
  enemies_number  : integer;
end record;
	function lfsr50(x : std_logic_vector(3 downto 0)) return std_logic_vector;
	function convSEG (N : std_logic_vector(3 downto 0)) return std_logic_vector;
	
end package;

package body NeonBlaster_pkg is
	function lfsr50(x : std_logic_vector(49 downto 0)) return std_logic_vector is
		begin
			return x(47 downto 0) & (x(0) xnor x(1) xnor x(4) xnor x(6)) & (x(8) xnor x(10) xnor x(13) xnor x(16));
		end function; 	
	function convSEG (N : std_logic_vector(3 downto 0)) return std_logic_vector is
		variable ans:std_logic_vector(6 downto 0);
begin
	Case N is
		when "0000" => ans:="1000000";	 
		when "0001" => ans:="1111001";
		when "0010" => ans:="0100100"; --
		when "0011" => ans:="0110000"; --
		when "0100" => ans:="0011001";
		when "0101" => ans:="0010010";
		when "0110" => ans:="0000010";
		when "0111" => ans:="1111000";
		when "1000" => ans:="0000000";
		when "1001" => ans:="0010000";	   
		when "1010" => ans:="0001000";
		when "1011" => ans:="0000011"; --
		when "1100" => ans:="1000110";
		when "1101" => ans:="0100001";
		when "1110" => ans:="0000110"; --
		when "1111" => ans:="0001110";				
		when others=> ans:="1111111";
	end case;	
	return ans;
end function convSEG;


end package body;